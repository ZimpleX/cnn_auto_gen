module addr_gen(clk,);
    parameter kern_buf_depth_addr = 16;

    reg 
endmodule
